`timescale 1ns / 1ps

// 실제로는 80Hz를 생성하는 코드
// 클럭 분주기 모듈 (Clock Divider)
// 방식: 카운터를 이용한 클럭 분주 (토글 방식)
module clock_8Hz(
    input i_clk,        
    input i_reset,
    output reg o_clk8Hz
    );

    // 카운터: 클럭 분주를 위한 카운터
    // 20비트로 선언 (2^20 = 1,048,576 > 625,000이므로 충분)
    reg [19:0] i_count=0;

    // 메인 로직: 클럭 상승엣지 또는 리셋 시 동작
    always @(posedge i_clk, posedge i_reset) begin
        // 비동기 리셋 처리
        if (i_reset) begin
            o_clk8Hz <= 0;
            i_count <= 0;
        end 
        
        // 정상 클럭 분주 동작
        else begin
            // 카운터가 목표값에 도달했는지 확인
            if (i_count == (1_250_000/2) - 1) begin // 8Hz : 12_500_000/2 = 6_250_000
                // 반주기 완료 -> 출력 클럭 토클 및 카운터 리셋
                i_count <= 0;
                o_clk8Hz <= ~o_clk8Hz;
            end 
            else begin
                // 아직 목표값 미달 -> 카운터 증가
                i_count <= i_count + 1;
            end
        end
    end
endmodule

    // =========================================================================
    // 클럭 분주 계산
    // =========================================================================
    // 목표: 100MHz → 8Hz 변환
    // 
    // 1) 8Hz 주기 계산:
    //    - 8Hz = 8 cycles/second
    //    - 한 주기 = 1/8 = 0.125초 = 125ms
    //    
    // 2) 100MHz에서 125ms에 해당하는 클럭 수:
    //    - 100,000,000 Hz × 0.125s = 12,500,000 클럭
    //    
    // 3) 토글 방식이므로 반주기마다 토글:
    //    - 12,500,000 ÷ 2 = 6,250,000 클럭마다 토글
    //    
    // 4) 카운터는 0부터 시작하므로:
    //    - 6,250,000 - 1 = 6,249,999까지 카운트
    // =========================================================================